ENTITY MouseHandlerTB IS
END MouseHandlerTB;

ARCHITECTURE TB OF MouseHandlerTB IS
BEGIN
